module p_encoder_32_5(in, out);

input 	[31:0] in;
output	[4:0] out;	 
// Because out being saved to in always_comb
logic 	[4:0] out;

always_comb begin

casex(in)

	32'b1:									begin out = 5'd0; end
	32'b1?:									begin out = 5'd1; end
	32'b1??:								begin out = 5'd2; end
	32'b1???:								begin out = 5'd3; end
	32'b1????:								begin out = 5'd4; end
	32'b1?????:								begin out = 5'd5; end
	32'b1??????:							begin out = 5'd6; end
	32'b1???????:							begin out = 5'd7; end
	32'b1????????:							begin out = 5'd8; end
	32'b1?????????:					 		begin out = 5'd9; end
	32'b1??????????:						begin out = 5'd10; end
	32'b1???????????:						begin out = 5'd11; end
	32'b1????????????:						begin out = 5'd12; end
	32'b1?????????????:						begin out = 5'd13; end
	32'b1??????????????:					begin out = 5'd14; end
	32'b1???????????????:					begin out = 5'd15; end
	32'b1????????????????:					begin out = 5'd16; end
	32'b1?????????????????:					begin out = 5'd17; end
	32'b1??????????????????:				begin out = 5'd18; end
	32'b1???????????????????:				begin out = 5'd19; end
	32'b1????????????????????:				begin out = 5'd20; end
	32'b1?????????????????????:				begin out = 5'd21; end
	32'b1??????????????????????:			begin out = 5'd22; end
	32'b1???????????????????????:			begin out = 5'd23; end
	32'b1????????????????????????:			begin out = 5'd24; end
	32'b1?????????????????????????:			begin out = 5'd25; end
	32'b1??????????????????????????:		begin out = 5'd26; end
	32'b1???????????????????????????:		begin out = 5'd27; end
	32'b1????????????????????????????:		begin out = 5'd28; end
	32'b1?????????????????????????????:		begin out = 5'd29; end
	32'b1??????????????????????????????:	begin out = 5'd30; end
	32'b1???????????????????????????????:	begin out = 5'd31; end
	default: out = 5'd0;
	endcase

end
endmodule

		