module p_encoder_32_5(in, out);

input 	[31:0] in;
output	[4:0] out;	 
// Because out being saved to in always_comb
logic 	[4:0] out;

always_comb begin

casex(in)

	32'b1:									begin out = 5'd0; end
	32'b1?:									begin out = 5'd1; end
	32'b1??:								begin out = 5'd2; end
	32'b1???:								begin out = 5'd3; end
	32'b1????:								begin out = 5'd4; end
	32'b1?????:								begin out = 5'd5; end
	32'b1??????:							begin out = 5'd6; end
	32'b1???????:							begin out = 5'd7; end
	32'b1????????:							begin out = 5'd8; end
	32'b1?????????:					 		begin out = 5'd9; end
	32'b1??????????:						begin out = 5'd10; end
	32'b1???????????:						begin out = 5'd11; end
	32'b1????????????:						begin out = 5'd12; end
	32'b1?????????????:						begin out = 5'd13; end
	32'b1??????????????:					begin out = 5'd14; end
	32'b1???????????????:					begin out = 5'd15; end
	32'b1????????????????:					begin out = 5'd16; end
	32'b1?????????????????:					begin out = 5'd17; end
	32'b1??????????????????:				begin out = 5'd18; end
	32'b1???????????????????:				begin out = 5'd19; end
	32'b1????????????????????:				begin out = 5'd20; end
	32'b1?????????????????????:				begin out = 5'd21; end
	32'b1??????????????????????:			begin out = 5'd22; end
	32'b1???????????????????????:			begin out = 5'd23; end
	32'b1????????????????????????:			begin out = 5'd24; end
	32'b1?????????????????????????:			begin out = 5'd25; end
	32'b1??????????????????????????:		begin out = 5'd26; end
	32'b1???????????????????????????:		begin out = 5'd27; end
	32'b1????????????????????????????:		begin out = 5'd28; end
	32'b1?????????????????????????????:		begin out = 5'd29; end
	32'b1??????????????????????????????:	begin out = 5'd30; end
	32'b1???????????????????????????????:	begin out = 5'd31; end
	default: out = 5'd0;
	endcase

end
endmodule

module decoder_5_32(in,out);

input 	[4:0] in;
output	[31:0] out;

logic [31:0] out;

always_comb begin

	if 		(in == 5'd0)	out = 32'b1;
	else if	(in == 5'd1)	out = 32'b10;
	else if (in == 5'd2)	out = 32'b100;
	else if (in == 5'd3)	out = 32'b1000;
	else if (in == 5'd4)	out = 32'b10000;
	else if (in == 5'd5)	out = 32'b100000;
	else if (in == 5'd6)	out = 32'b1000000;
	else if (in == 5'd7)	out = 32'b10000000;
	else if (in == 5'd8)	out = 32'b100000000;
	else if (in == 5'd9)	out = 32'b1000000000;
	else if (in == 5'd10)	out = 32'b10000000000;
	else if (in == 5'd11)	out = 32'b100000000000;
	else if (in == 5'd12)	out = 32'b1000000000000;
	else if (in == 5'd13)	out = 32'b10000000000000;
	else if (in == 5'd14)	out = 32'b100000000000000;
	else if (in == 5'd15)	out = 32'b1000000000000000;
	else if (in == 5'd16)	out = 32'b10000000000000000;
	else if (in == 5'd17)	out = 32'b100000000000000000;
	else if (in == 5'd18)	out = 32'b1000000000000000000;
	else if (in == 5'd19)	out = 32'b10000000000000000000;
	else if (in == 5'd20)	out = 32'b100000000000000000000;
	else if (in == 5'd21)	out = 32'b1000000000000000000000;
	else if (in == 5'd22)	out = 32'b10000000000000000000000;
	else if (in == 5'd23)	out = 32'b100000000000000000000000;
	else if (in == 5'd24)	out = 32'b1000000000000000000000000;
	else if (in == 5'd25)	out = 32'b10000000000000000000000000;
	else if (in == 5'd26)	out = 32'b100000000000000000000000000;
	else if (in == 5'd27)	out = 32'b1000000000000000000000000000;
	else if (in == 5'd28)	out = 32'b10000000000000000000000000000;
	else if (in == 5'd29)	out = 32'b100000000000000000000000000000;
	else if (in == 5'd30)	out = 32'b1000000000000000000000000000000;
	else if (in == 5'd31)	out = 32'b10000000000000000000000000000000;

end
endmodule

module one_hot_32(in,out);

input [31:0] in;
wire [4:0] out1;
output [31:0] out;

p_encoder_32_5 enc1 (in,out1);
decoder_5_32   dec1 (out1,out);

endmodule

module scientific(in, mantissa, exponent);

input 	[31:0] in;
output	[7:0] mantissa;
output	[4:0] exponent;

logic 	[4:0] exponent;
logic 	[31:0] hot_out, and_result, exponent_bits, hot_copy;
logic 	[7:0] mantissa;
logic 	bit_test;

one_hot_32 hot1 (in,hot_out);	

always_comb 
begin
	hot_copy = hot_out;

	if ( hot_copy >= 32'd128) 
	begin
		for( int i = 7; i >= 0; i--) 
			begin 
			and_result = in & hot_copy;
			mantissa[i] = |and_result;
			hot_copy = hot_copy >> 1;
			end
			//hot_copy = hot_copy << 1; Why didn't this work?

			hot_copy = hot_copy << 1;
	end
		
	else 
	begin
		mantissa = in;
		hot_copy = 32'd0;
	end

end

p_encoder_32_5 exponent_enc(hot_copy,exponent);	

endmodule
		
